// Based on https://github.com/B-Lang-org/bsc-contrib Copyright (c) 2020 Bluespec, Inc. All rights reserved.
// SPDX-License-Identifier: BSD-3-Clause
// Modified by Kamyar Mohajerani

package Bus;

import BusDefines :: *;
import BusFIFO    :: *;

export BusDefines :: *;
export BusFIFO    :: *;

endpackage
