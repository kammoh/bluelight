package SIPO;

import Vector::*;
import PISO::*;

export SIPO::*;
export Vector::*;

interface SIPO #(numeric type size, type el_type);
  method Action enq(el_type in_data); 
  method Action deq;
  (* always_ready *)
  method CountType#(size) count;
  (* always_ready *)
  method Bool isFull;
  (* always_ready *)
  method Bool notFull;
  (* always_ready *)
  method Vector#(size, el_type) data;
endinterface

// Pipelined SIPO (Serial In, Parallel Out)
// if full enq can happen simultanously with deq of first element 
module mkPipelineSIPO (SIPO#(size, el_type)) provisos (Bits#(el_type, el_type_sz));
  Reg#(Vector#(size, el_type)) vec <- mkRegU;
  Reg#(CountType#(size)) count_reg <- mkReg(0);
  RWire#(el_type) rwEnq <- mkRWire();
  let pwDeq <- mkPulseWire();

  Bool full = count_reg == fromInteger(valueOf(size));
  
  (* fire_when_enabled, no_implicit_conditions *)
  rule update if (isValid(rwEnq.wget) || pwDeq);
    case (rwEnq.wget) matches
      tagged Valid .v:
        begin
          vec <= shiftInAtN(vec, v);
          if (pwDeq) // simultanous enq & deq
            count_reg <= 1;
          else // enq only
            count_reg <= count_reg + 1;
        end
      tagged Invalid: // deq only
        count_reg <= 0;
    endcase
  endrule

  method Action enq(el_type el) if (!full || pwDeq);
    rwEnq.wset(el);
  endmethod
        
  method Action deq if (full);
    pwDeq.send();
  endmethod

  method Vector#(size, el_type) data;
    return vec;
  endmethod

  method CountType#(size) count;
    return count_reg;
  endmethod

  method Bool isFull;
    return full;
  endmethod

  method Bool notFull;
    return !full;
  endmethod
endmodule : mkPipelineSIPO


module mkSIPO (SIPO#(size, el_type)) provisos (Bits#(el_type, el_type_sz));
  Reg#(Vector#(size, el_type)) vec <- mkRegU;
  Reg#(CountType#(size)) count_reg <- mkReg(0);

  Bool full = count_reg == fromInteger(valueOf(size));

  method Action enq(el_type v) if (!full);
    vec <= shiftInAtN(vec, v);
    count_reg <= count_reg + 1;
  endmethod
        
  method Action deq if (full);
    count_reg <= 0;
  endmethod

  method Vector#(size, el_type) data;
    return vec;
  endmethod

  method CountType#(size) count;
    return count_reg;
  endmethod

  method Bool isFull;
    return full;
  endmethod

  method Bool notFull;
    return !full;
  endmethod

endmodule : mkSIPO



interface MyShiftReg #(numeric type size, type el_type);
  (* always_ready *)
  method Action enq(el_type in_data); 
  (* always_ready *)
  method Vector#(size, el_type) data;
endinterface

module mkMyShiftReg (MyShiftReg#(size, el_type)) provisos (Bits#(el_type, el_type_sz));
  Reg#(Vector#(size, el_type)) vec <- mkRegU;

  method Action enq(el_type v);
    vec <= shiftInAtN(vec, v);
  endmethod
  method Vector#(size, el_type) data;
    return vec;
  endmethod
endmodule : mkMyShiftReg

endpackage : SIPO