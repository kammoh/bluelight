package Bus;

import BusDefines :: *;
import BusFIFO    :: *;


export BusDefines :: *;
export BusFIFO    :: *;

endpackage
